../chisel/verilog/register_template.v